
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity ROM_Memory is

  Port ( 
         ADDRESS : in STD_LOGIC_VECTOR (7 downto 0);
         DATA : out STD_LOGIC_VECTOR (31 downto 0);
         ENABLE : in STD_LOGIC;
         CLK : in STD_LOGIC);

end ROM_Memory;


architecture Behavioral of ROM_Memory is 


type myTab_type is array( 0 to 255) of std_logic_vector(31 downto 0);
signal romfile  :   myTab_type;


begin 

	romfile(0) <= "00000000000000000000000000000110";
	romfile(1) <= "01000000000000000000000000010001";
	romfile(2) <= "10000000000000000000000000000000";
	romfile(3) <= "10000000000000000000000000000000";
	romfile(4) <= "10000000000000000000000000000000";
	romfile(5) <= "10000000000000000000000000000000";
	romfile(6) <= "10000000000000000000000000000000";
	romfile(7) <= "10000000000000000000000000000000";
	romfile(8) <= "10000000000000000000000000000000";
	romfile(9) <= "10000000000000000000000000000000";
	romfile(10) <= "10000000000000000000000000000000";
	romfile(11) <= "10000000000000000000000000000000";
	romfile(12) <= "10000000000000000000000000000000";
	romfile(13) <= "10000000000000000000000000000000";
	romfile(14) <= "10000000000000000000000000000000";
	romfile(15) <= "10000000000000000000000000000000";
	romfile(16) <= "10000000000000000000000000000000";
	romfile(17) <= "10000000000000000000000000000000";
	romfile(18) <= "10000000000000000000000000000000";
	romfile(19) <= "10000000000000000000000000000000";
	romfile(20) <= "10000000000000000000000000000000";
	romfile(21) <= "10000000000000000000000000000000";
	romfile(22) <= "10000000000000000000000000000000";
	romfile(23) <= "10000000000000000000000000000000";
	romfile(24) <= "10000000000000000000000000000000";
	romfile(25) <= "10000000000000000000000000000000";
	romfile(26) <= "10000000000000000000000000000000";
	romfile(27) <= "10000000000000000000000000000000";
	romfile(28) <= "10000000000000000000000000000000";
	romfile(29) <= "10000000000000000000000000000000";
	romfile(30) <= "10000000000000000000000000000000";
	romfile(31) <= "10000000000000000000000000000000";
	romfile(32) <= "10000000000000000000000000000000";
	romfile(33) <= "10000000000000000000000000000000";	
	romfile(34) <= "10000000000000000000000000000000";
	romfile(35) <= "10000000000000000000000000000000";
	romfile(36) <= "10000000000000000000000000000000";
	romfile(37) <= "10000000000000000000000000000000";
	romfile(38) <= "10000000000000000000000000000000";
	romfile(39) <= "10000000000000000000000000000000";
	romfile(40) <= "10000000000000000000000000000000";
	romfile(41) <= "10000000000000000000000000000000";
	romfile(42) <= "10000000000000000000000000000000";
	romfile(43) <= "10000000000000000000000000000000";
	romfile(44) <= "10000000000000000000000000000000";
	romfile(45) <= "10000000000000000000000000000000";
	romfile(46) <= "10000000000000000000000000000000";
	romfile(47) <= "10000000000000000000000000000000";
	romfile(48) <= "10000000000000000000000000000000";
	romfile(49) <= "10000000000000000000000000000000";
	romfile(50) <= "10000000000000000000000000000000";
	romfile(51) <= "10000000000000000000000000000000";
	romfile(52) <= "10000000000000000000000000000000";
	romfile(53) <= "10000000000000000000000000000000";
	romfile(54) <= "10000000000000000000000000000000";
	romfile(55) <= "10000000000000000000000000000000";
	romfile(56) <= "10000000000000000000000000000000";
	romfile(57) <= "10000000000000000000000000000000";
	romfile(58) <= "10000000000000000000000000000000";
	romfile(59) <= "10000000000000000000000000000000";
	romfile(60) <= "10000000000000000000000000000000";
	romfile(61) <= "10000000000000000000000000000000";
	romfile(62) <= "10000000000000000000000000000000";
	romfile(63) <= "10000000000000000000000000000000";
	romfile(64) <= "10000000000000000000000000000000";
	romfile(65) <= "10000000000000000000000000000000";
	romfile(66) <= "10000000000000000000000000000000";
	romfile(67) <= "10000000000000000000000000000000";
	romfile(68) <= "10000000000000000000000000000000";
	romfile(69) <= "10000000000000000000000000000000";
	romfile(70) <= "10000000000000000000000000000000";
	romfile(71) <= "10000000000000000000000000000000";
	romfile(72) <= "10000000000000000000000000000000";
	romfile(73) <= "10000000000000000000000000000000";
	romfile(74) <= "10000000000000000000000000000000";
	romfile(75) <= "10000000000000000000000000000000";
	romfile(76) <= "10000000000000000000000000000000";
	romfile(77) <= "10000000000000000000000000000000";
	romfile(78) <= "10000000000000000000000000000000";
	romfile(79) <= "10000000000000000000000000000000";
	romfile(80) <= "10000000000000000000000000000000";
	romfile(81) <= "10000000000000000000000000000000";
	romfile(82) <= "10000000000000000000000000000000";
	romfile(83) <= "10000000000000000000000000000000";
	romfile(84) <= "10000000000000000000000000000000";
	romfile(85) <= "10000000000000000000000000000000";
	romfile(86) <= "10000000000000000000000000000000";
	romfile(87) <= "10000000000000000000000000000000";
	romfile(88) <= "10000000000000000000000000000000";
	romfile(89) <= "10000000000000000000000000000000";
	romfile(90) <= "10000000000000000000000000000000";
	romfile(91) <= "10000000000000000000000000000000";
	romfile(92) <= "10000000000000000000000000000000";
	romfile(93) <= "10000000000000000000000000000000";
	romfile(94) <= "10000000000000000000000000000000";
	romfile(95) <= "10000000000000000000000000000000";
	romfile(96) <= "10000000000000000000000000000000";
	romfile(97) <= "10000000000000000000000000000000";
	romfile(98) <= "10000000000000000000000000000000";
	romfile(99) <= "10000000000000000000000000000000";
	romfile(100) <= "10000000000000000000000000000000";
	romfile(101) <= "10000000000000000000000000000000";
	romfile(102) <= "10000000000000000000000000000000";
	romfile(103) <= "10000000000000000000000000000000";
	romfile(104) <= "10000000000000000000000000000000";
	romfile(105) <= "10000000000000000000000000000000";
	romfile(106) <= "10000000000000000000000000000000";
	romfile(107) <= "10000000000000000000000000000000";
	romfile(108) <= "10000000000000000000000000000000";
	romfile(109) <= "10000000000000000000000000000000";
	romfile(110) <= "10000000000000000000000000000000";
	romfile(111) <= "10000000000000000000000000000000";
	romfile(112) <= "10000000000000000000000000000000";
	romfile(113) <= "10000000000000000000000000000000";
	romfile(114) <= "10000000000000000000000000000000";
	romfile(115) <= "10000000000000000000000000000000";
	romfile(116) <= "10000000000000000000000000000000";
	romfile(117) <= "10000000000000000000000000000000";
	romfile(118) <= "10000000000000000000000000000000";
	romfile(119) <= "10000000000000000000000000000000";
	romfile(120) <= "10000000000000000000000000000000";
	romfile(121) <= "10000000000000000000000000000000";
	romfile(122) <= "10000000000000000000000000000000";
	romfile(123) <= "10000000000000000000000000000000";
	romfile(124) <= "10000000000000000000000000000000";
	romfile(125) <= "10000000000000000000000000000000";
	romfile(126) <= "10000000000000000000000000000000";
	romfile(127) <= "10000000000000000000000000000000";
	romfile(128) <= "10000000000000000000000000000000";
	romfile(129) <= "10000000000000000000000000000000";
	romfile(130) <= "10000000000000000000000000000000";
	romfile(131) <= "10000000000000000000000000000000";
	romfile(132) <= "10000000000000000000000000000000";
	romfile(133) <= "10000000000000000000000000000000";
	romfile(134) <= "10000000000000000000000000000000";
	romfile(135) <= "10000000000000000000000000000000";
	romfile(136) <= "10000000000000000000000000000000";
	romfile(137) <= "10000000000000000000000000000000";
	romfile(138) <= "10000000000000000000000000000000";
	romfile(139) <= "10000000000000000000000000000000";
	romfile(140) <= "10000000000000000000000000000000";
	romfile(141) <= "10000000000000000000000000000000";
	romfile(142) <= "10000000000000000000000000000000";
	romfile(143) <= "10000000000000000000000000000000";
	romfile(144) <= "10000000000000000000000000000000";
	romfile(145) <= "10000000000000000000000000000000";
	romfile(146) <= "10000000000000000000000000000000";
	romfile(147) <= "10000000000000000000000000000000";
	romfile(148) <= "10000000000000000000000000000000";
	romfile(149) <= "10000000000000000000000000000000";
	romfile(150) <= "10000000000000000000000000000000";
	romfile(151) <= "10000000000000000000000000000000";
	romfile(152) <= "10000000000000000000000000000000";
	romfile(153) <= "10000000000000000000000000000000";
	romfile(154) <= "10000000000000000000000000000000";
	romfile(155) <= "10000000000000000000000000000000";
	romfile(156) <= "10000000000000000000000000000000";
	romfile(157) <= "10000000000000000000000000000000";
	romfile(158) <= "10000000000000000000000000000000";
	romfile(159) <= "10000000000000000000000000000000";
	romfile(160) <= "10000000000000000000000000000000";
	romfile(161) <= "10000000000000000000000000000000";
	romfile(162) <= "10000000000000000000000000000000";
	romfile(163) <= "10000000000000000000000000000000";
	romfile(164) <= "10000000000000000000000000000000";
	romfile(165) <= "10000000000000000000000000000000";
	romfile(166) <= "10000000000000000000000000000000";
	romfile(167) <= "10000000000000000000000000000000";
	romfile(168) <= "10000000000000000000000000000000";
	romfile(169) <= "10000000000000000000000000000000";
	romfile(170) <= "10000000000000000000000000000000";
	romfile(171) <= "10000000000000000000000000000000";
	romfile(172) <= "10000000000000000000000000000000";
	romfile(173) <= "10000000000000000000000000000000";
	romfile(174) <= "10000000000000000000000000000000";
	romfile(175) <= "10000000000000000000000000000000";
	romfile(176) <= "10000000000000000000000000000000";
	romfile(177) <= "10000000000000000000000000000000";
	romfile(178) <= "10000000000000000000000000000000";
	romfile(179) <= "10000000000000000000000000000000";
	romfile(180) <= "10000000000000000000000000000000";
	romfile(181) <= "10000000000000000000000000000000";
	romfile(182) <= "10000000000000000000000000000000";
	romfile(183) <= "10000000000000000000000000000000";
	romfile(184) <= "10000000000000000000000000000000";
	romfile(185) <= "10000000000000000000000000000000";
	romfile(186) <= "10000000000000000000000000000000";
	romfile(187) <= "10000000000000000000000000000000";
	romfile(188) <= "10000000000000000000000000000000";
	romfile(189) <= "10000000000000000000000000000000";
	romfile(190) <= "10000000000000000000000000000000";
	romfile(191) <= "10000000000000000000000000000000";
	romfile(192) <= "10000000000000000000000000000000";
	romfile(193) <= "10000000000000000000000000000000";
	romfile(194) <= "10000000000000000000000000000000";
	romfile(195) <= "10000000000000000000000000000000";
	romfile(196) <= "10000000000000000000000000000000";
	romfile(197) <= "10000000000000000000000000000000";
	romfile(198) <= "10000000000000000000000000000000";
	romfile(199) <= "10000000000000000000000000000000";
	romfile(200) <= "10000000000000000000000000000000";
	romfile(201) <= "10000000000000000000000000000000";
	romfile(202) <= "10000000000000000000000000000000";
	romfile(203) <= "10000000000000000000000000000000";
	romfile(204) <= "10000000000000000000000000000000";
	romfile(205) <= "10000000000000000000000000000000";
	romfile(206) <= "10000000000000000000000000000000";
	romfile(207) <= "10000000000000000000000000000000";
	romfile(208) <= "10000000000000000000000000000000";
	romfile(209) <= "10000000000000000000000000000000";
	romfile(210) <= "10000000000000000000000000000000";
	romfile(211) <= "10000000000000000000000000000000";
	romfile(212) <= "10000000000000000000000000000000";
	romfile(213) <= "10000000000000000000000000000000";
	romfile(214) <= "10000000000000000000000000000000";
	romfile(215) <= "10000000000000000000000000000000";
	romfile(216) <= "10000000000000000000000000000000";
	romfile(217) <= "10000000000000000000000000000000";
	romfile(218) <= "10000000000000000000000000000000";
	romfile(219) <= "10000000000000000000000000000000";
	romfile(220) <= "10000000000000000000000000000000";
	romfile(221) <= "10000000000000000000000000000000";
	romfile(222) <= "10000000000000000000000000000000";
	romfile(223) <= "10000000000000000000000000000000";
	romfile(224) <= "10000000000000000000000000000000";
	romfile(225) <= "10000000000000000000000000000000";
	romfile(226) <= "10000000000000000000000000000000";
	romfile(227) <= "10000000000000000000000000000000";
	romfile(228) <= "10000000000000000000000000000000";
	romfile(229) <= "10000000000000000000000000000000";
	romfile(230) <= "10000000000000000000000000000000";
	romfile(231) <= "10000000000000000000000000000000";
	romfile(232) <= "10000000000000000000000000000000";
	romfile(233) <= "10000000000000000000000000000000";
	romfile(234) <= "10000000000000000000000000000000";
	romfile(235) <= "10000000000000000000000000000000";
	romfile(236) <= "10000000000000000000000000000000";
	romfile(237) <= "10000000000000000000000000000000";
	romfile(238) <= "10000000000000000000000000000000";
	romfile(239) <= "10000000000000000000000000000000";
	romfile(240) <= "10000000000000000000000000000000";
	romfile(241) <= "10000000000000000000000000000000";
	romfile(242) <= "10000000000000000000000000000000";
	romfile(243) <= "10000000000000000000000000000000";
	romfile(244) <= "10000000000000000000000000000000";
	romfile(245) <= "10000000000000000000000000000000";
	romfile(246) <= "10000000000000000000000000000000";
	romfile(247) <= "10000000000000000000000000000000";
	romfile(248) <= "10000000000000000000000000000000";
	romfile(249) <= "10000000000000000000000000000000";
	romfile(250) <= "10000000000000000000000000000000";
	romfile(251) <= "10000000000000000000000000000000";
	romfile(252) <= "10000000000000000000000000000000";
	romfile(253) <= "10000000000000000000000000000000";
	romfile(254) <= "10000000000000000000000000000000";
	romfile(255) <= "10000000000000000000000000000000";

    react: Process (enable, clk) is

    begin

    -- if (enable = '0') then

          -- enable action here
	  -- ???????

     if rising_edge(clk) then

          -- clock edge reaction here

            DATA <= romfile(to_integer(unsigned(ADDRESS)));
          
      end if;

   
    end process react;


end Behavioral;


