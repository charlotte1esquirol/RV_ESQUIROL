library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;



entity byte_extend is



  Port (Din :  in STD_LOGIC_VECTOR (7 downto 0);
    	Dout : out STD_LOGIC_VECTOR (31 downto 0);
	unsigned1 : in STD_LOGIC);       


end byte_extend;

architecture Behavioral of byte_extend is



alias MSB : std_logic is Din ( 7 );
alias sigsize : std_logic_vector is Dout ( 7 downto 0 );
alias sigzero : std_logic_vector is Dout ( 31 downto 8 );


begin

	process ( Din, unsigned1 )

	begin

	if ( unsigned1 = '1' or MSB = '0' ) then

		sigzero <= "000000000000000000000000";
		sigsize <= Din;


	else 
		sigzero <= "111111111111111111111111"; 
		sigsize <= Din;


	end if;

	end process;
		

end Behavioral;

