library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity StateMachine_tb is

end StateMachine_tb; 


architecture Behavioral of StateMachine_tb is

component StateMachine

	port
	(
		clk : in std_logic;
		rst	 : in	std_logic;
		trigger	 : in	std_logic;
		PREADY	 : in	std_logic;
		unaligned : in std_logic;
		op1 : out std_logic;
		op2 : out std_logic;
		first_cycle : out std_logic;
		busy_sel : out std_logic_vector (1 downto 0) ;
		preq_sel : out std_logic;
		PENABLE : out std_logic);

end component; 

     


signal sbusy : STD_LOGIC_VECTOR(1 downto 0);

signal sCLK, sRST, strigger, sPREADY, sunaligned, sop1, sop2, sfirst, sPENABLE, spreq : STD_LOGIC; 



begin 



UUT : StateMachine port map ( clk=>sCLK, rst=>sRST, trigger=>strigger, PREADY=>sPREADY, unaligned=>sunaligned, op1=>sop1, op2=>sop2, first_cycle=>sfirst, preq_sel=>spreq, busy_sel=>sbusy, PENABLE => sPENABLE );



process 

    begin

    sCLK <='0';

        wait for 10 ns;

    sCLK <='1';

        wait for 10 ns;

    end process;





process

    begin 

    -- on commence par un reset pour tout bien mettre � 0

	sRST<='1';
	wait for 30 ns;

    -- cas o� on reste � s0

   	sRST<='0'; 

	strigger<='0';

        sPREADY<='0';

        sunaligned<='0';
        
        wait for 30 ns;

     -- cas o� on passe � s1 et y reste

        strigger<='1';

        wait for 30 ns; 

     -- cas o� on revient � s1 et repasse � s0 au prochain clock edge

        sPREADY<='1'; 

        wait for 40 ns; 

     -- cas o� on passe � s2 et ensuite forcement � s3 puis � s0

        sunaligned<='1';

        wait for 200 ns;

     end process;

end Behavioral;

        








