library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
use work.rv_esquirol_pkg.all;

-- prototype defined in 'neorv32_package.vhd'
package rv_esquirol_controlunit_image_pkg is

constant control_unit_image : mem32_t := (

x"00000006",
x"40000011",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000",
x"80000000");

end rv_esquirol_controlunit_image_pkg;
